module f_sub(
	input [1599:0] absorb_outcome,
	input [7:0] rc,
	output [1599:0] s_out
);
integer i,j,k;



reg [63:0] a [24:0];
reg [63:0] b [4:0];
reg [63:0] d [4:0];
reg [63:0] e [24:0];

reg [63:0] a1 [24:0];

reg [1599:0] out;

wire [63:0] rc_wire;

/*************************************************
*   Name :          rc_wire
*   Description:    transfer 8bits ROUND CONSTANTS into 64 bits ROUND CONSTANTS
*************************************************/

assign rc_wire={rc[7],31'b0,rc[6],15'b0,rc[5],7'b0,rc[4],3'b0,rc[3:0]}; 

always @(*) begin

/*************************************************
*   Name :          a
*   Description:    assign absorb_outcome to a from 0 bit to 1599 bit，every a[i] is 64 bits
*************************************************/

	for(i=0;i<25;i=i+1)
		a[i]=absorb_outcome[((i<<6))+:64]; 

/*************************************************
*   Name :          b
*   Description:    assign (j,0) xor (j,1) xor (j,2) xor (j,3) xor (j,4) to b[j]，every b[j] is 64 bits (Theta first step)
*************************************************/

	for(j=0;j<5;j=j+1)
		b[j]=a[j]^a[5+j]^a[10+j]^a[15+j]^a[20+j];

/*************************************************
*   Name :          d
*   Description:    assign b[(x-1) mod 5, z] xor b[(x+1) mod 5, (z-1) mod 64] to d[i]，every d[i] is 64 bits (Theta second step)
*************************************************/ 

	d[0]=b[4]^{b[1][62:0],b[1][63]};
	d[1]=b[0]^{b[2][62:0],b[2][63]};
	d[2]=b[1]^{b[3][62:0],b[3][63]};
	d[3]=b[2]^{b[4][62:0],b[4][63]};
	d[4]=b[3]^{b[0][62:0],b[0][63]};

/*************************************************
*   Name :          a1
*   Description:    assign Theta second step to a1[i]，every a[i] is 64 bits
*************************************************/

	a1[0]=a[0]^d[0];

/*************************************************
*   Name :          b
*   Description:    assign Rho & Pi to b[i]，every b[i] is 64 bits 
*************************************************/

	b[0]=a1[0];
	a1[6]=a[6]^d[1];
	b[1]={a1[6][19:0],a1[6][63:20]};
	a1[12]=a[12]^d[2];
	b[2]={a1[12][20:0],a1[12][63:21]};
	a1[18]=a[18]^d[3];
	b[3]={a1[18][42:0],a1[18][63:43]};
	a1[24]=a[24]^d[4];
	b[4]={a1[24][49:0],a1[24][63:50]};

/*************************************************
*   Name :          e
*   Description:    assign Chi & Iota to e[i]，every e[i] is 64 bits
*************************************************/

	e[0]=b[0]^((~b[1]) & b[2]);
	e[0]=e[0]^rc_wire;
	e[1]=b[1]^((~b[2]) & b[3]);
	e[2]=b[2]^((~b[3]) & b[4]);
	e[3]=b[3]^((~b[4]) & b[0]);
	e[4]=b[4]^((~b[0]) & b[1]);


	a1[3]=a[3]^d[3];
	b[0]={a1[3][35:0],a1[3][63:36]};
	a1[9]=a[9]^d[4];
	b[1]={a1[9][43:0],a1[9][63:44]};
	a1[10]=a[10]^d[0];
	b[2]={a1[10][60:0],a1[10][63:61]};
	a1[16]=a[16]^d[1];
	b[3]={a1[16][18:0],a1[16][63:19]};
	a1[22]=a[22]^d[2];
	b[4]={a1[22][2:0],a1[22][63:3]};
	e[5]=b[0]^((~b[1]) & b[2]);
	e[6]=b[1]^((~b[2]) & b[3]);
	e[7]=b[2]^((~b[3]) & b[4]);
	e[8]=b[3]^((~b[4]) & b[0]);
	e[9]=b[4]^((~b[0]) & b[1]);



	a1[1]=a[1]^d[1];
	b[0]={a1[1][62:0],a1[1][63]};
	a1[7]=a[7]^d[2];
	b[1]={a1[7][57:0],a1[7][63:58]};
	a1[13]=a[13]^d[3];
	b[2]={a1[13][38:0],a1[13][63:39]};
	a1[19]=a[19]^d[4];
	b[3]={a1[19][55:0],a1[19][63:56]};
	a1[20]=a[20]^d[0];
	b[4]={a1[20][45:0],a1[20][63:46]};
	e[10]=b[0]^((~b[1]) & b[2]);
	e[11]=b[1]^((~b[2]) & b[3]);
	e[12]=b[2]^((~b[3]) & b[4]);
	e[13]=b[3]^((~b[4]) & b[0]);
	e[14]=b[4]^((~b[0]) & b[1]);


	a1[4]=a[4]^d[4];
	b[0]={a1[4][36:0],a1[4][63:37]};
	a1[5]=a[5]^d[0];
	b[1]={a1[5][27:0],a1[5][63:28]};
	a1[11]=a[11]^d[1];
	b[2]={a1[11][53:0],a1[11][63:54]};
	a1[17]=a[17]^d[2];
	b[3]={a1[17][48:0],a1[17][63:49]};
	a1[23]=a[23]^d[3];
	b[4]={a1[23][7:0],a1[23][63:8]};
	e[15]=b[0]^((~b[1]) & b[2]);
	e[16]=b[1]^((~b[2]) & b[3]);
	e[17]=b[2]^((~b[3]) & b[4]);
	e[18]=b[3]^((~b[4]) & b[0]);
	e[19]=b[4]^((~b[0]) & b[1]);


	a1[2]=a[2]^d[2];
	b[0]={a1[2][1:0],a1[2][63:2]};
	a1[8]=a[8]^d[3];
	b[1]={a1[8][8:0],a1[8][63:9]};
	a1[14]=a[14]^d[4];
	b[2]={a1[14][24:0],a1[14][63:25]};
	a1[15]=a[15]^d[0];
	b[3]={a1[15][22:0],a1[15][63:23]};
	a1[21]=a[21]^d[1];
	b[4]={a1[21][61:0],a1[21][63:62]};
	e[20]=b[0]^((~b[1]) & b[2]);
	e[21]=b[1]^((~b[2]) & b[3]);
	e[22]=b[2]^((~b[3]) & b[4]);
	e[23]=b[3]^((~b[4]) & b[0]);
	e[24]=b[4]^((~b[0]) & b[1]);

/*************************************************
*   Name :          out
*   Description:    assign e[0]~e[24] to out from 0 bit to 1599 bit
*************************************************/

	for(i=0;i<25;i=i+1)
		out[((i<<6))+:64]=e[i];

end

/*************************************************
*   Name :          s_out
*   Description:    assign out to s_out
*************************************************/

assign s_out=out;


endmodule